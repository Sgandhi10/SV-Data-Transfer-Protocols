/******************************************************************************
* Filename : I2C_Peripheral.sv
* Author : Soham Gandhi
* Date : 1/17/2025
* Description : This file contains the I2C Peripheral(Slave) module.
* Version : 1.0 (SG) Initial Version
******************************************************************************/

module I2C_Peripheral(
    
)