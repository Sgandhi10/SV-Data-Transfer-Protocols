/*******************************************************************************
* File: 8b10b_encoder.sv
* Author: Soham Gandhi
* Date: 2025-08-03
* Description: This is a 8b10b encoder known for being used in high speed communication.
*   This converter will be implemented based on the spec mentioned here: 
* Version: 1.0
*******************************************************************************/

module 8b10b_encoder #() (
    input   logic       clk,
    input   logic       rst_n,

    input   logic [7:0] data_in,
    output  logic [7:0] data_out
);

// 

endmodule