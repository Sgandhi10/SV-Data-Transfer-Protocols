/*******************************************************************************
* File: 8b10b_decoder.sv
* Author: Soham Gandhi
* Date: 2025-08-03
* Description:
* Version: 1.0
*******************************************************************************/

